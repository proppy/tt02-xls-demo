module user_module(
  input wire [7:0] io_in,
  output wire [7:0] io_out
);
  assign io_out = io_in;
endmodule
